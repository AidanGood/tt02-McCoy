/*
* Aidan Good
* alu.v
* The ALU. Only operation is addition currently.
*/

module alu(
	input [5:0] op1,
	input [5:0] op2,
	output [5:0] aluOut);
    
    assign aluOut = op1 + op2;
	

	
endmodule


